`timescale 1ns/10ps
`include "./src/struct_s.sv"
`include "./src/stats_reg.sv"



